library verilog;
use verilog.vl_types.all;
entity UART_tb is
end UART_tb;
